library verilog;
use verilog.vl_types.all;
entity Datapath_tb is
end Datapath_tb;
